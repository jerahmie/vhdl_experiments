library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity clk_1 is
  port ( clk_in : in STD_LOGIC;
	reset  : in STD_LOGIC;
	clk_out : out STD_LOGIC );
end clk_1;
architecture Behavioral of clk_1 is
  signal temporal : STD_LOGIC;
  signal counter : integer range 0 to 124999 := 0;
begin  -- Behavioral of clk_1
  frequency_divider: process (reset, clk_in)
  begin
    if reset = '1' then
      temporal <= '0';
      counter <= 0;
    elsif rising_edge(clk_in) then
      if counter = 10 then
        temporal <= NOT(temporal);
        counter <= 0;
        else
          counter <= counter + 1;
      end if;
    end if;
  end process;
  
  clk_out <= temporal;
end Behavioral;
